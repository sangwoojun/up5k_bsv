typedef Bit#(32) Word;
typedef Bit#(5) RIndx;
typedef Bit#(3) SizeType;

